`define  NONE       
`define  MODE_64     
`define  NONE       
`define  NONE       
`define  VCS       
`define  SIM       
`define  NONE       
`define  NONE       
`define  NONE       
`define  NONE       
`define  TILE_MODEL 
`define  SFU_MODEL 
`define  VIT_LUT 
